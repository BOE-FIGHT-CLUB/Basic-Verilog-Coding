//========================================
//
//  Verilog Tamplate Module
//
// sync with https://github.com/BigKuchz/Basic-Verilog-Coding.git
//
//
//========================================

module boe_fight_club_top(

);



endmodule