//========================================
//
//  Verilog Tamplate Module
//
//========================================

module boe_fight_club_top(

);

endmodule